module data_memory(
	input clk,
	input w_en,
	input [3:0] addr,
	input [3:0] data_in,
	output [3:0] data_out);
	
endmodule
