module program_sequencer(
	//IO
	);
	
endmodule
