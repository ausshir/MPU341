library verilog;
use verilog.vl_types.all;
entity test_instruction_decoder is
end test_instruction_decoder;
