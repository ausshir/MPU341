module data_memory(
	//IO
	);
	
endmodule
