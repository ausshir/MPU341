library verilog;
use verilog.vl_types.all;
entity test_bench_for_instruction_decoder is
end test_bench_for_instruction_decoder;
