module computational_unit(
	//IO
	);
	
endmodule
