library verilog;
use verilog.vl_types.all;
entity test_program_memory is
end test_program_memory;
