library verilog;
use verilog.vl_types.all;
entity test_program_sequencer is
end test_program_sequencer;
