library verilog;
use verilog.vl_types.all;
entity test_program_sequencer_2 is
end test_program_sequencer_2;
